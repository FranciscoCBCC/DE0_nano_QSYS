LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY DE0_NANO IS
	PORT ( 
		CLOCK_50 : IN STD_LOGIC);
END DE0_NANO;

ARCHITECTURE arch OF DE0_NANO IS
BEGIN

	PROCESS(CLOCK_50)
		BEGIN

		END PROCESS;

END arch;